magic
tech scmos
timestamp 788836334
<< nwell >>
rect 43 104 157 210
rect 19 11 181 83
<< pdiffusion >>
rect 42 56 43 64
rect 42 55 90 56
rect 42 39 46 55
rect 49 51 79 52
rect 49 43 50 51
rect 78 43 79 51
rect 49 42 79 43
rect 82 39 90 55
rect 42 36 90 39
rect 42 28 43 36
rect 110 59 166 60
rect 118 37 119 59
rect 122 52 154 56
rect 122 44 126 52
rect 150 44 154 52
rect 122 40 154 44
rect 157 37 158 59
rect 110 36 166 37
rect 132 28 146 36
<< metal1 >>
rect 7 48 8 77
rect 3 46 8 48
rect 0 0 8 8
rect 16 86 17 94
rect 30 72 31 80
rect 42 65 43 68
rect 42 64 90 65
rect 42 56 43 64
rect 94 68 106 109
rect 183 86 184 94
rect 169 72 170 80
rect 94 60 110 68
rect 94 59 166 60
rect 42 36 45 56
rect 94 52 110 59
rect 49 51 110 52
rect 49 43 50 51
rect 78 43 110 51
rect 49 42 110 43
rect 42 28 43 36
rect 30 16 31 24
rect 22 15 94 16
rect 16 0 17 8
rect 98 0 102 42
rect 118 55 158 59
rect 118 41 123 55
rect 118 37 132 41
rect 110 36 132 37
rect 135 24 143 44
rect 153 41 158 55
rect 146 37 158 41
rect 146 36 166 37
rect 170 24 178 25
rect 106 15 178 16
rect 183 0 184 8
rect 192 49 193 78
rect 192 0 200 8
<< metal2 >>
rect 0 78 200 80
rect 0 77 193 78
rect 0 48 3 77
rect 7 69 193 77
rect 7 65 43 69
rect 90 65 193 69
rect 7 49 193 65
rect 197 49 200 78
rect 7 48 200 49
rect 0 46 200 48
rect 42 37 86 46
rect 0 15 200 33
rect 0 11 20 15
rect 94 11 106 15
rect 178 11 200 15
rect 0 0 200 11
<< pdcontact >>
rect 34 28 42 68
rect 43 56 90 64
rect 50 43 78 51
rect 43 28 90 36
rect 110 60 166 68
rect 110 37 118 59
rect 126 44 150 52
rect 158 37 166 59
rect 110 28 132 36
rect 146 28 166 36
<< m2contact >>
rect 3 48 7 77
rect 43 65 90 69
rect 20 11 94 15
rect 106 11 178 15
rect 193 49 197 78
<< psubstratepcontact >>
rect 8 0 16 94
rect 17 86 89 94
rect 111 86 183 94
rect 17 0 93 8
rect 107 0 183 8
rect 184 0 192 94
<< nsubstratencontact >>
rect 22 16 30 80
rect 31 72 90 80
rect 110 72 169 80
rect 31 16 94 24
rect 170 25 178 80
rect 106 16 178 24
<< psubstratepdiff >>
rect 0 0 8 8
rect 16 86 17 94
rect 89 86 111 94
rect 183 86 184 94
rect 16 0 17 8
rect 93 0 107 8
rect 183 0 184 8
rect 192 0 200 8
<< nsubstratendiff >>
rect 30 72 31 80
rect 90 72 110 80
rect 169 72 170 80
rect 30 16 31 24
rect 94 16 106 72
rect 170 24 178 25
<< pad >>
rect 50 109 150 209
<< labels >>
rlabel space 0 0 200 210 1 mbb
rlabel metal2 4 15 4 15 3 Vdd
rlabel m2contact 3 56 3 56 3 GND
<< end >>
