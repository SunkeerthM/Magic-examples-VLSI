magic
tech scmos
timestamp 1625909441
<< nwell >>
rect -4 -1 17 20
<< polysilicon >>
rect 5 11 8 13
rect 5 -4 8 2
rect 7 -8 8 -4
rect 5 -17 8 -8
rect 5 -29 8 -27
<< ndiffusion >>
rect 2 -21 5 -17
rect -2 -27 5 -21
rect 8 -21 10 -17
rect 14 -21 17 -17
rect 8 -27 17 -21
<< pdiffusion >>
rect -1 7 5 11
rect 3 3 5 7
rect -1 2 5 3
rect 8 8 15 11
rect 8 4 10 8
rect 14 4 15 8
rect 8 2 15 4
<< metal1 >>
rect 3 15 11 19
rect -1 7 3 15
rect 10 -4 14 4
rect -6 -8 3 -4
rect 10 -8 22 -4
rect 10 -17 14 -8
rect -2 -32 2 -21
rect 2 -36 9 -32
rect 13 -36 18 -32
<< ntransistor >>
rect 5 -27 8 -17
<< ptransistor >>
rect 5 2 8 11
<< polycontact >>
rect 3 -8 7 -4
<< ndcontact >>
rect -2 -21 2 -17
rect 10 -21 14 -17
<< pdcontact >>
rect -1 3 3 7
rect 10 4 14 8
<< psubstratepcontact >>
rect -2 -36 2 -32
rect 9 -36 13 -32
rect 18 -36 22 -32
<< nsubstratencontact >>
rect -1 15 3 19
rect 11 15 15 19
<< labels >>
rlabel metal1 7 17 7 17 5 Vdd
rlabel metal1 0 -6 0 -6 3 a
rlabel metal1 16 -6 16 -6 1 b
rlabel metal1 6 -34 6 -34 1 gnd
<< end >>
